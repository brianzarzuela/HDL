-- Brian Zarzuela
-- Lab 5

entity gen_add_sub is
end gen_add_sub;